module top_module (
    input a,
    input b,
    input c,
    input d,
    output q 
);
    

endmodule

// bd
// dc
// bcd
// ad
// ac
// acd
// abd
// abc
// abcd
